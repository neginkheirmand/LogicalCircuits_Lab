`timescale 1ns / 1ps
module decoder4to16TestBench;
	reg [3:0] in;
	reg en;
	wire [15:0] dout;
	Decoder4to16 uut (
		.in(in), 
		.en(en), 
		.dout(dout)
	);
	initial begin
	//enable 1
	en = 1'b1;
	//0 0 0 0 
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b0;
		#100;
	//0 0 0 1
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b1;
		#100;
	//0 0 1 0
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b1;
	in[3]=1'b0;
		#100;
	//0 0 1 1
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b1;
	in[3]=1'b1;
		#100;
	//0 1 0 0
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b0;
	in[3]=1'b0;
		#100;
	//0 1 0 1
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b0;
	in[3]=1'b1;
		#100;
	//0 1 1 0
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b1;
	in[3]=1'b0;
		#100;
	//0 1 1 1
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b1;
	in[3]=1'b1;
		#100;
	//1 0 0 0 
	in[0]=1'b1;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b0;
		#100;
	//1 0 0 1
	in[0]=1'b1;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b1;

		#100;
	//enable 0
	en = 1'b0;
	//0 0 0 0 
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b0;
		#100;
	//0 0 0 1
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b1;
		#100;
	//0 0 1 0
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b1;
	in[3]=1'b0;
		#100;
	//0 0 1 1
	in[0]=1'b0;
	in[1]=1'b0;
	in[2]=1'b1;
	in[3]=1'b1;
		#100;
	//0 1 0 0
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b0;
	in[3]=1'b0;
		#100;
	//0 1 0 1
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b0;
	in[3]=1'b1;
		#100;
	//0 1 1 0
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b1;
	in[3]=1'b0;
		#100;
	//0 1 1 1
	in[0]=1'b0;
	in[1]=1'b1;
	in[2]=1'b1;
	in[3]=1'b1;
		#100;
	//1 0 0 0 
	in[0]=1'b1;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b0;
		#100;
	//1 0 0 1
	in[0]=1'b1;
	in[1]=1'b0;
	in[2]=1'b0;
	in[3]=1'b1;
		#100;
      

	end
      
endmodule

