`timescale 1ns / 1ps
module PriorityModuleTestbBench;
	reg D3;
	reg D2;
	reg D1;
	reg D0;
	wire A1;
	wire A0;
	MyPriorityEncoder uut (
		.D3(D3), 
		.D2(D2), 
		.D1(D1), 
		.D0(D0), 
		.A1(A1), 
		.A0(A0)
	);
	initial begin
	//0 0 0 0 
		D3 = 1'b0; D2 = 1'b0; D1 = 1'b0; D0 = 1'b0;
		#100;
	//0 0 0 1
		D3 = 1'b0; D2 = 1'b0; D1 = 1'b0; D0 = 1'b1;
		#100;
	//0 0 1 0 
		D3 = 1'b0; D2 = 1'b0; D1 = 1'b1; D0 = 1'b0;
		#100;
	//0 0 1 1 
		D3 = 1'b0; D2 = 1'b0; D1 = 1'b1; D0 = 1'b1;
		#100;
	//0 1 0 0 
		D3 = 1'b0; D2 = 1'b1; D1 = 1'b0; D0 = 1'b0;
		#100;
	//0 1 0 1 
		D3 = 1'b0; D2 = 1'b1; D1 = 1'b0; D0 = 1'b1;
		#100;
	//0 1 1 0 
		D3 = 1'b0; D2 = 1'b1; D1 = 1'b1; D0 = 1'b0;
		#100;
	//0 1 1 1 
		D3 = 1'b0; D2 = 1'b1; D1 = 1'b1; D0 = 1'b1;
		#100;
	//1 0 0 0 
		D3 = 1'b1; D2 = 1'b0; D1 = 1'b0; D0 = 1'b0;
		#100;
	//1 0 0 1 
		D3 = 1'b1; D2 = 1'b0; D1 = 1'b0; D0 = 1'b1;
		#100;
	//1 0 1 0 
		D3 = 1'b1; D2 = 1'b0; D1 = 1'b1; D0 = 1'b0;
		#100;
	//1 0 1 1 
		D3 = 1'b1; D2 = 1'b0; D1 = 1'b1; D0 = 1'b1;
		#100;
	//1 1 0 0 
		D3 = 1'b1; D2 = 1'b1; D1 = 1'b0; D0 = 1'b0;
		#100;
	//1 1 0 1 
		D3 = 1'b1; D2 = 1'b1; D1 = 1'b0; D0 = 1'b1;
		#100;
	//1 1 1 0 
		D3 = 1'b1; D2 = 1'b1; D1 = 1'b1; D0 = 1'b0;
		#100;
	//1 1 1 1 
		D3 = 1'b1; D2 = 1'b1; D1 = 1'b1; D0 = 1'b1;
		#100;

		$finish;
	end
      
endmodule

