`timescale 1ns / 1ps
module SequenceDetectorTestBench(
    );


endmodule
